`timescale 1ns/100ps
module flopr_tb;
    
    int counter, errors;
    logic clk, rst;
    integer file;
    
	logic clock, reset, d, q, q_esperado;
    
    parameter max_vectors = 19;
    logic [30:0] vectors[max_vectors];

    flopr dut(clock, reset, d, q);

    initial begin
        counter = 0; errors = 0;
		rst = 1'b1; #12; rst = 0;
		clk=0;
		
		if(~rst) begin
			$readmemb("flopr.tv", vectors);
		end	
		
		file = $fopen("flopr_out.txt");
    
        $display("Iniciando Testbench");
        $display("---------------");
        $display("| Clk | Rst | d | q |");
        
        $fwrite(file, "Iniciando Testbench\n");
        $fwrite(file, "---------------\n");
        $fwrite(file, "| Clk | Rst | d | q |\n"); 	
    end
	        
    always begin
        clk = 1; #6;
        clk = 0; #5;
    end

    always @(posedge clk) begin
        if(~rst) begin
	        {clock, reset, d, q_esperado} = vectors[counter];
        end
	end

    always @(negedge clk)	//Sempre (que o clock descer)
        if(~rst) begin
			if(q_esperado !== 1'bx) begin

				assert (q === q_esperado) begin
					$display("|  %b  |  %b  | %b | %b | OK", clock, reset, d, q);
					$fwrite(file, "|  %b  |  %b  | %b | %b | OK\n", clock, reset, d, q);
				end else begin
					//Mostra mensagem de erro se a saída do DUT for diferente da saída esperada
					$error("q = %b (%b esperado) {Linha %d}", q, q_esperado, counter+1);
								
					errors = errors + 1; //Incrementa contador de erros a cada bit errado encontrado
				end
	
				if(counter+1 == max_vectors) begin
					$display("Testes Efetuados  = %0d", counter+1);
					$display("Erros Encontrados = %0d", errors);
					$fwrite(file, "Testes Efetuados  = %0d\n", counter+1);
					$fwrite(file, "Erros Encontrados = %0d\n", errors);
					#10
					$stop;
				end    
			end
			counter++; //Incrementa contador dos vertores de teste
        end
endmodule
 
 
