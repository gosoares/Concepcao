`timescale 1ns/100ps
module adder_tb;
    
    int counter, errors, aux_error;
    logic clk, rst;
    integer file;
    
    logic a, b, cin, s, s_esperado, cout, cout_esperado;
    
    parameter max_vectors = 8;
    logic [4:0] vectors[max_vectors];

    adder dut(a, b, cin, s, cout);

    initial begin
        counter = 0; errors = 0;
		rst = 1'b1; #12; rst = 0;
		clk=0;
		
		if(~rst) begin
			$readmemb("adder.tv", vectors);
		end	
		
		file = $fopen("adder_out.txt");
    
        $display("Iniciando Testbench");
        $display("---------------");
        $display("| A | B | Cin | S |");
        
        $fwrite(file, "Iniciando Testbench");
        $fwrite(file, "---------------");
        $fwrite(file, "| A | B | Cin | S |"); 	
    end
	        
    always begin
        clk = 1; #7;
        clk = 0; #5;
    end

    always @(posedge clk)
        if(~rst) begin
	        {a, b, cin, cout_esperado, s_esperado} = vectors[counter];	
        end

    always @(negedge clk)	//Sempre (que o clock descer)
        if(~rst && s_esperado !== 1'bx && cout_esperado !== 1'bx) begin
            aux_error = errors;
            
            assert (s === s_esperado) else begin
                errors++;
                $error("| %b | %b |  %b  | %b |  %b  | ERROR: S = %b", a, b, cin, s_esperado, cout_esperado, s);
                $fwrite(file, "| %b | %b |  %b  | %b |  %b  | ERROR: S = %b", a, b, cin, s_esperado, cout_esperado, s);
            end
            
            assert (s === s_esperado) else begin
                errors++;
                $error("| %b | %b |  %b  | %b |  %b  | ERROR: Cout = %b", a, b, cin, s_esperado, cout_esperado, cout);
                $fwrite(file, "| %b | %b |  %b  | %b |  %b  | ERROR: Cout = %b", a, b, cin, s_esperado, cout_esperado, cout);
            end

            if(aux_error === errors) begin // Nao houve erro
                $display("| %b | %b |  %b  | %b |  %b  | OK", a, b, cin, s, cout);
                $fwrite(file, "| %b | %b |  %b  | %b |  %b  | OK", a, b, cin, s, cout);
            end

            counter++;	//Incrementa contador dos vertores de teste
            if(counter == max_vectors) begin
	            $display("Testes Efetuados  = %0d", counter);
	            $display("Erros Encontrados = %0d", errors);
	            $fwrite(file, "Testes Efetuados  = %0d", counter);
	            $fwrite(file, "Erros Encontrados = %0d", errors);
	            #10
	            $stop;
            end     
        end
endmodule
 
 
